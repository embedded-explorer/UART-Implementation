//----------------------------------------------------------------------------
// Title       : Micro UART Controller
// Design      : UART Receiver
// File        : uart_rx.sv
//----------------------------------------------------------------------------
// Description : UART Receiver module, responsible to receive incoming serial 
//               data on RX line and write 8 bit parallel data to RX FIFO
//----------------------------------------------------------------------------
// Author      :
// Version     : 1.0 - Initial Version
//               2.0 - Added subset of control and status features from 16550
//                     Renamed and restructured FIFO write logic for convinience
//----------------------------------------------------------------------------

`timescale 1ns/1ns

module uart_rx(
  // Clock and reset
  input                 uart_clk_i        , // reference input clock
  input                 uart_rst_n_i      , // active low synchronous reset
  input                 rx_clk_en_i       , // RX clock enable pulse 16 times baud rate

  // Data output to RX FIFO
  output  logic  [9:0]  rx_fifo_data_o    , // RX FIFO data bus
  output  logic         rx_fifo_wr_en_o   , // RX FIFO write enable
  
  // Control and status signals
  input          [1:0]  word_len_i        , // Number Data Bits
  input                 parity_en_i       , // Parity Enable
  input                 even_parity_sel_i , // Select even parity
  input                 stp_bits_i        , // Number of stop bits
  output  logic         rsr_full_o        , // RX shift register is filled
    
  // Serial data input
  input                 uart_rx_i           // UART RX input Pin
);

//----------------------------------------------------------------------------
// Custom data types
//----------------------------------------------------------------------------
  
  // FSM State Encoding
  typedef enum logic [4:0]{
    S_IDLE   = 5'b00001,
    S_START  = 5'b00010,
    S_DATA   = 5'b00100,
    S_PARITY = 5'b01000,
    S_STOP   = 5'b10000
  } state_coding_t;

  state_coding_t curr_state ; // FSM current state register
  state_coding_t next_state ; // FSM next state register

//----------------------------------------------------------------------------
// Internal signal decleration
//----------------------------------------------------------------------------

  logic [2:0] bit_count       ; // counter to count number of bits received
  logic [3:0] tik_count       ; // counter to count number of rx enable ticks
  logic [7:0] data            ; // receiver shift register
  logic [7:0] data_rcvd       ; // Data received, to be written to FIFO
  logic       check_bit       ; // calculated check bit - even parity
  logic       parity_rcvd     ; // received parity
  logic       parity_err      ; // parity error detected
  logic       frame_err       ; // Frame error detected
  logic       stop_bit_1_done ; // Flag used to stay in stop state
  logic       rx_fifo_wr_en   ; // Enable writing to RX FIFO
  logic       rx_fifo_wr_en_d ; // delay write enable signal by 1 cycle
  
  // Signals used for clock synchronization  
  logic       uart_rx_d0      ;
  logic       uart_rx_d1      ;
  logic       uart_rx_d2      ;
  
//----------------------------------------------------------------------------
// Combinational Logic
//----------------------------------------------------------------------------
  
  // Wriet enable generated by fifo write logic will be high for 1/16 baud period
  // read enable given to FIFO must be high only for 1 clock cycle
  // detect positive edge on write enable to make it high for only one cycle
  assign rx_fifo_wr_en_o = (rx_fifo_wr_en & !rx_fifo_wr_en_d);
  
  // Assign data received based on the word length selected
  assign data_rcvd = (word_len_i == 2'b11) ? data : data[7:1];
  
  // Parity error detection logic
  always_comb begin
    if(parity_en_i) begin
    // When parity is enabled
      if(even_parity_sel_i) begin
      // When even parity is selected
        if(check_bit) begin
        // When received parity and calculated check bit are not equal
          parity_err = 1'b1; // parity error is generated
        end else begin
          parity_err = 1'b0;
        end
      end else begin
      // When odd parity is selected
        if(check_bit) begin
          parity_err = 1'b0;
        end else begin
        // When received parity and calculated check bit are not equal
          parity_err = 1'b1; // parity error is generated
        end
      end
    end else begin
      parity_err = 1'b0;
    end
  end
  
  // Frame error detection logic
  always_ff @(posedge uart_clk_i)begin
    if(!uart_rst_n_i) begin
      frame_err <= 1'b0 ;
    end else begin
      if((curr_state == S_STOP) && (tik_count == 4'hE)) begin
      // Check for frame error in stop state at center of baud interval
        if(!uart_rx_d2) begin
        // If rx line is low this indicates invalid stop bit
          frame_err <= 1'b1; // frame error is detected
        end else begin
          frame_err <= 1'b0 ;
        end
      end else begin
        frame_err <= 1'b0 ;
      end
    end
  end
  
//----------------------------------------------------------------------------
// Sequential Logic
//----------------------------------------------------------------------------
  
  // As UART is asynchronous received data will not synchronized to reference clock
  // hence synchronize the received data to reference clock
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
      uart_rx_d0 <= 1'b0;
      uart_rx_d1 <= 1'b0;
      uart_rx_d2 <= 1'b0;
    end else begin
      if(rx_clk_en_i) begin
        uart_rx_d0 <= uart_rx_i ;
        uart_rx_d1 <= uart_rx_d0;
        uart_rx_d2 <= uart_rx_d1;
      end
    end
  end
  
  // Check bit calculation for parity
  always_ff @(posedge uart_clk_i)begin
    if (!uart_rst_n_i) begin
      check_bit <= 1'b0;
    end else begin
      if(curr_state == S_STOP) begin
      // Calculate check bit for parity
        check_bit <= parity_rcvd ^ (data_rcvd);
      end
    end
  end
    
  // FIFO write logic
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
    // Clear signals on reset
      rx_fifo_wr_en  <= 1'b0  ;
      rx_fifo_data_o <= 10'h0 ;
    end else begin
      if((curr_state == S_STOP) && (tik_count == 4'hF)) begin
      // Check whether center of baud interval is reached in stop state
      // received data along with parity error and frame error is written
        rx_fifo_data_o  <= {frame_err, parity_err, data_rcvd};
        if(stp_bits_i) begin
        // In 2 stop bit mode
          if(stop_bit_1_done) begin
          // Data is written to RX FIFO after receiving 2 stop bits
            rx_fifo_wr_en <= 10'h1 ;
          end else begin
            rx_fifo_wr_en <= 10'h0 ;
          end
        end else begin
        // In 1 stop bit mode data is written after 1 stop bit
          rx_fifo_wr_en <= 10'h1 ;
        end
      end else begin
        rx_fifo_data_o <= 10'h0 ;
        rx_fifo_wr_en  <= 10'h0 ;
      end
    end
  end
  
  // Delay write enable pulse by 1 cycle to detect edge of write enable
  always_ff @(posedge uart_clk_i)begin
    if (!uart_rst_n_i) begin
      rx_fifo_wr_en_d <= 1'b0;
    end else begin
      rx_fifo_wr_en_d <= rx_fifo_wr_en;
    end
  end
    
//----------------------------------------------------------------------------
// Finite State Machine
//----------------------------------------------------------------------------
  
  // Sequential Present state logic
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
      curr_state <= S_IDLE    ; // Upon reset move to IDLE state
    end else begin
      curr_state <= next_state; // Synchronously change the state
    end
  end
  
  // Combinational next state decoder
  always_comb begin
    if(rx_clk_en_i) begin
    // Sample rx line only on reception of tx clock enable pulse
      case(curr_state)
      // Next state will be decided by checking current state
            
        S_IDLE  : begin
          if (uart_rx_d2 & !uart_rx_d1) begin
          // Dettect falling edge on rx line
            next_state = S_START ; // move to start state
          end else begin
          // Wait in IDLE state until start bit is detected on RX line
            next_state = S_IDLE  ;
          end
        end
            
        S_START : begin
          if (tik_count >= 4'h6) begin
          // Check whether center of baud interval is reached
            if (!uart_rx_d2) begin
            // check start at center of baud interval
              next_state = S_DATA ; // move to DATA state, if rx is still low
            end else begin
            // If start bit is high, indicates invalid start bit
              next_state = S_IDLE ; // move to IDLE state
            end
          end else begin
          // Wait until center of baud interval is reached
            next_state = S_START ; // move to START state
          end
        end
            
        S_DATA  : begin
          if ((bit_count >= (word_len_i + 4)) && (tik_count >= 4'hF)) begin
          // Check whether complete word is received and center of baud interval is reached
            if(parity_en_i) begin
            // When parity is enabled
              next_state = S_PARITY ; // move to PARITY state
            end else begin
            // When parity is not enabled
              next_state = S_STOP   ; // move to STOP state
            end
          end else begin
          // stay in data state until comple word is received
            next_state = S_DATA ;
          end
        end
                
        S_PARITY : begin
          if (tik_count >= 4'hF) begin
          // Wait until center of baud interval is reached
            next_state = S_STOP  ; // move to STOP state
          end else begin
          // Stay is parity state until center of baud interval is reached
            next_state = S_PARITY;
          end
        end
                
        S_STOP  : begin
          if(tik_count >= 4'hF) begin
          // When center of baud interval is reached
            if (stp_bits_i & !stop_bit_1_done) begin
            // When 2 stop bit mode is selected and first stop bit is not transmitted
              next_state = S_STOP ; // stay in stop state for 1 more interval
            end else begin
            // When all stop bits are transmitted
              next_state = S_IDLE ; // move to idle state
            end
          end else begin
          // Stay in stop state until center of baud interval is reached
            next_state = S_STOP ;
          end
        end
                
        default : next_state = S_IDLE ;
                
      endcase
    end else begin
      next_state = curr_state  ; // Stay in present state
    end
  end
  
  // Sequential output and register logic
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
    // Clear the signals on reset
      bit_count       <= 3'b0 ;
      tik_count       <= 4'h0 ;
      data            <= 8'h0 ;
      parity_rcvd     <= 1'b0 ;
      stop_bit_1_done <= 1'b0 ;
      rsr_full_o      <= 1'b0 ;
    end else begin
      if (rx_clk_en_i) begin
      // When receiver clcok enable is high
        case(curr_state)
        
          S_IDLE  : begin
          // Clear the signals in idle state
            bit_count       <= 3'b0 ;
            data            <= 8'h0 ;
            parity_rcvd     <= 1'b0 ;
            stop_bit_1_done <= 1'b0 ;
            rsr_full_o      <= 1'b0 ;
          end
          
          S_START : begin
            if (tik_count >= 4'h6) begin
            // When RX tick count is reached to 7
              tik_count      <= 4'h0 ; // clear tick count
            end else begin
            // When RX tick count is not yet reached to 7
              tik_count <= tik_count + 1'b1 ; // increment tick count
            end
          end

          S_DATA  : begin         
            if (tik_count >= 4'hF) begin
            // When RX tick count is reached 15 
            // sample incoming RX data at center of baud interval
              tik_count <= 1'b0                    ; // clear tick count
              data      <= {uart_rx_d2, data[7:1]} ; // shift incoming data bit into receiver shift register
              bit_count <= bit_count + 1'b1        ; // increment bit count on receiving each bit
            end else begin
            // If TX tick count is not yet reached to 15
              tik_count <= tik_count + 1'b1 ; // increment tick count
            end
          end
          
          S_PARITY :begin
            bit_count <= 3'b0             ; // Clear bit count
            if (tik_count >= 4'hF) begin
            // Sample parity bit at center of baud interval
              parity_rcvd <= uart_rx_d2;
              tik_count   <= 4'h0      ;
            end else begin
              tik_count   <= tik_count + 1'b1 ; // Increment tick count
            end
          end
          
          S_STOP  : begin
            rsr_full_o      <= 1'b1 ; // Indicate RX shift register is filled
            tik_count       <= tik_count + 1'b1 ; // Increment tick count
            if (tik_count >= 4'hE) begin
              stop_bit_1_done <= 1'b1 ; // Indicate stop state is entered
            end
          end
          
        endcase
      end
    end
  end

endmodule