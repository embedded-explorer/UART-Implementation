//----------------------------------------------------------------------------
// Title       : Micro UART Controller
// Design      : UART Transmitter
// File        : uart_tx.sv
//----------------------------------------------------------------------------
// Description : UART transmitter module, responsible to read parallel data 
//               from TX FIFO and shift out bits serailly over TX line
//----------------------------------------------------------------------------
// Author      :
// Version     : 1.0 - Initial Version
//               2.0 - Added subset of control and status features from 16550
//                     Renamed few signals for convinience
//----------------------------------------------------------------------------

`timescale 1ns/1ns

module uart_tx(
  // Clock and reset
  input                 uart_clk_i        , // reference input clock
  input                 uart_rst_n_i      , // active low synchronous reset
  input                 tx_clk_en_i       , // TX clock enable pulse at baud rate

  // Data input from TX FIFO
  input          [7:0]  tx_fifo_data_i    , // TX FIFO data bus
  input                 tx_fifo_empty_i   , // TX FIFO empty
  output  logic         tx_fifo_rd_en_o   , // TX FIFO read enable
  
  // Control and status signals
  input          [1:0]  word_len_i        , // Number Data Bits
  input                 parity_en_i       , // Parity Enable
  input                 even_parity_sel_i , // Select even parity
  input                 stp_bits_i        , // Number of stop bits
  output  logic         tsr_empty_o       , // TX Shift register empty
  
  // Serial data output
  output  logic         uart_tx_o           // UART TX output Pin
);

//----------------------------------------------------------------------------
// Custom data types
//----------------------------------------------------------------------------

  // FSM State Encoding
  typedef enum logic [4:0]{
    S_IDLE   = 5'b00001,
    S_START  = 5'b00010,
    S_DATA   = 5'b00100,
    S_PARITY = 5'b01000,
    S_STOP   = 5'b10000
  } state_coding_t;

  state_coding_t curr_state ; // FSM current state register
  state_coding_t next_state ; // FSM next state register

//----------------------------------------------------------------------------
// Internal signal decleration
//----------------------------------------------------------------------------

  logic [2:0] bit_count       ; // counter to count number of bits shifted
  logic [7:0] data            ; // internal transmit shift register
  logic       tx_fifo_rd_en   ; // enable to read data from tx fifo
  logic       tx_fifo_rd_en_d ; // delay read enable signal by 1 cycle
  logic       check_bit       ; // calculated parity check bit
  logic       parity_bit      ; // parity calulated locally
  logic       stop_bit_1_done ; // Flag used to stay in stop state
  
//----------------------------------------------------------------------------
// Combinational Logic
//----------------------------------------------------------------------------

  // Read enable generated by FSM will be high for 1 baud period
  // read enable given to FIFO must be high only for 1 clock cycle
  // detect positive edge on read enable to make it high for only one cycle
  assign tx_fifo_rd_en_o = (tx_fifo_rd_en & !tx_fifo_rd_en_d);
  
  // Transmit shift register is empty when tx is in idle state
  assign tsr_empty_o = (curr_state == S_IDLE) ? 1'b1 : 1'b0;

//----------------------------------------------------------------------------
// Sequential Logic
//----------------------------------------------------------------------------

  // Delay read enable pulse by 1 cycle to detect edge of write enable
  always_ff @(posedge uart_clk_i)begin
    if (!uart_rst_n_i) begin
      tx_fifo_rd_en_d <= 1'b0;
    end else begin
      tx_fifo_rd_en_d <= tx_fifo_rd_en;
    end
  end
  
  // Check bit calculation for parity
  always_ff @(posedge uart_clk_i)begin
    if (!uart_rst_n_i) begin
      check_bit <= 1'b0;
    end else begin
      if (tx_fifo_rd_en_o) begin
        case(word_len_i)
        // Calculate check bit for parity
        // Number of bits on which parity is calculated depends on number of data bits
          2'b10   : check_bit <= ^tx_fifo_data_i[6:0]; // 7-Data bits
          2'b11   : check_bit <= ^tx_fifo_data_i     ; // 8-Data bits
          default : check_bit <= 1'b0;
        endcase
      end
    end
  end
  
  // Parity generation based on selection
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
      parity_bit <= 1'b0;
    end else begin
      if(even_parity_sel_i) begin
      // Even parity must be generated
        parity_bit <= check_bit;
      end else begin
      // Odd parity must be generated
        parity_bit <= ~check_bit;
      end
    end
  end
  
//----------------------------------------------------------------------------
// Finite State Machine
//----------------------------------------------------------------------------

  // Sequential Present state logic
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
      curr_state <= S_IDLE    ; // Upon reset move to IDLE state
    end else begin
      curr_state <= next_state; // Synchronously change the state
    end
  end

  // Combinational next state decoder
  always_comb begin
    if(tx_clk_en_i) begin
    // Enable transmission only on reception of tx clock enable pulse
      case(curr_state)
      // Next state will be decided by checking current state
      
        S_IDLE  : begin
          if (!tx_fifo_empty_i) begin
          // When data is avilable in TX FIFO
            next_state = S_START ; // move to START state
          end else begin
          // When TX FIFO is empty
            next_state = S_IDLE  ; // Stay in IDLE state
          end
        end
        
        S_START : begin
          next_state = S_DATA ; // move to DATA state unconditionally
        end
        
        S_DATA  : begin
          if (bit_count >= (word_len_i + 4)) begin
          // on sending out complete word
            if(parity_en_i) begin
            // Check whether parity is enabled
              next_state = S_PARITY ; // move to PARITY state
            end else begin
              next_state = S_STOP   ; // move to STOP state
            end
          end else begin
          // Stay in data state until comple word is transmitted
            next_state = S_DATA ;
          end
        end
        
        S_PARITY : begin
          next_state = S_STOP ; // move to STOP state
        end
        
        S_STOP  : begin
          if(stp_bits_i & !stop_bit_1_done) begin
          // When 2 stop bit mode is selected and first stop bit is not transmitted
            next_state = S_STOP; // stay in stop state for 1 more cycle
          end else begin
            if (!tx_fifo_empty_i) begin
            // When data is avilable in TX FIFO
              next_state = S_START ; // move to START state
            end else begin
            // When TX FIFO is empty
              next_state = S_IDLE  ; // move to IDLE state
            end
          end
        end
        
        default : next_state = S_IDLE  ;
        
      endcase
    end else begin
      next_state = curr_state  ; // Stay in present state
    end
  end

  // Sequential output and register logic
  always_ff @(posedge uart_clk_i) begin
    if (!uart_rst_n_i) begin
    // Clear the signals on reset
      bit_count       <= 3'b0 ;
      data            <= 1'b0 ;
      tx_fifo_rd_en   <= 1'b0 ;
      uart_tx_o       <= 1'b1 ;
      stop_bit_1_done <= 1'b0 ;
    end else begin
      if (tx_clk_en_i) begin
      // signals will be changed only when tx clock enable pulse is present
        case(curr_state)
        // Output signals will be based on the current state
        
          S_IDLE  : begin
            uart_tx_o       <= 1'b1 ; // TX line is held high during IDLE state
            stop_bit_1_done <= 1'b0 ;
          end
          
          S_START : begin
            stop_bit_1_done <= 1'b0           ;
            uart_tx_o       <= 1'b0           ; // send start bit (high to low)
            tx_fifo_rd_en   <= 1'b1           ; // generate read enable signal
            data            <= tx_fifo_data_i ; // load data read from FIFO to transmit shift register
          end
          
          S_DATA  : begin
            tx_fifo_rd_en <= 1'b0            ; // clear read enable
            uart_tx_o     <= data[bit_count] ; // send out bit indexed by bit count
            bit_count     <= bit_count + 1'b1; // increment bit count on sending each bit
          end
          
          S_PARITY :begin
            bit_count <= 1'b0      ; // bit count is cleared
            uart_tx_o <= parity_bit; // Transmit parity bit
            // Uncomment below line for parity checking
            //uart_tx_o <= 1'b0      ; // Transmit wrong parity bit
          end
          
          S_STOP  : begin
            stop_bit_1_done <= 1'b1   ; // Indicate first stop bit is transmitted
            bit_count       <= 3'h0   ; // bit count is cleared
            uart_tx_o       <= 1'b1   ; // send stop bit (x to high)
            // Uncomment below line for testing frame error
            //uart_tx_o       <= 1'b0   ; // send invalid stop bit
          end

        endcase
      end
    end
  end

endmodule